
module ProjectFile (
	clk_clk,
	regs_export,
	reset_reset_n);	

	input		clk_clk;
	output	[7:0]	regs_export;
	input		reset_reset_n;
endmodule
