// ProjectFile.v

// Generated using ACDS version 20.1 720

`timescale 1 ps / 1 ps
module ProjectFile (
		input  wire       alarm_active_switch_export, // alarm_active_switch.export
		input  wire       clk_clk,                    //                 clk.clk
		input  wire       down_button_export,         //         down_button.export
		input  wire       edit_alarm_switch_export,   //   edit_alarm_switch.export
		input  wire       edit_time_switch_export,    //    edit_time_switch.export
		input  wire       edit_timer_switch_export,   //   edit_timer_switch.export
		output wire [9:0] leds_export,                //                leds.export
		input  wire       left_button_export,         //         left_button.export
		input  wire       reset_reset_n,              //               reset.reset_n
		input  wire       right_button_export,        //        right_button.export
		input  wire       save_switch_export,         //         save_switch.export
		output wire [7:0] segment1_export,            //            segment1.export
		output wire [7:0] segment2_export,            //            segment2.export
		output wire [7:0] segment3_export,            //            segment3.export
		output wire [7:0] segment4_export,            //            segment4.export
		output wire [7:0] segment5_export,            //            segment5.export
		output wire [7:0] segment6_export,            //            segment6.export
		input  wire       timer_active_switch_export, // timer_active_switch.export
		input  wire       uart_rxd,                   //                uart.rxd
		output wire       uart_txd,                   //                    .txd
		input  wire       up_button_export            //           up_button.export
	);

	wire  [31:0] cpu_data_master_readdata;                             // mm_interconnect_0:CPU_data_master_readdata -> CPU:d_readdata
	wire         cpu_data_master_waitrequest;                          // mm_interconnect_0:CPU_data_master_waitrequest -> CPU:d_waitrequest
	wire         cpu_data_master_debugaccess;                          // CPU:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:CPU_data_master_debugaccess
	wire  [15:0] cpu_data_master_address;                              // CPU:d_address -> mm_interconnect_0:CPU_data_master_address
	wire   [3:0] cpu_data_master_byteenable;                           // CPU:d_byteenable -> mm_interconnect_0:CPU_data_master_byteenable
	wire         cpu_data_master_read;                                 // CPU:d_read -> mm_interconnect_0:CPU_data_master_read
	wire         cpu_data_master_write;                                // CPU:d_write -> mm_interconnect_0:CPU_data_master_write
	wire  [31:0] cpu_data_master_writedata;                            // CPU:d_writedata -> mm_interconnect_0:CPU_data_master_writedata
	wire  [31:0] cpu_instruction_master_readdata;                      // mm_interconnect_0:CPU_instruction_master_readdata -> CPU:i_readdata
	wire         cpu_instruction_master_waitrequest;                   // mm_interconnect_0:CPU_instruction_master_waitrequest -> CPU:i_waitrequest
	wire  [15:0] cpu_instruction_master_address;                       // CPU:i_address -> mm_interconnect_0:CPU_instruction_master_address
	wire         cpu_instruction_master_read;                          // CPU:i_read -> mm_interconnect_0:CPU_instruction_master_read
	wire         mm_interconnect_0_jtag_avalon_jtag_slave_chipselect;  // mm_interconnect_0:JTAG_avalon_jtag_slave_chipselect -> JTAG:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_avalon_jtag_slave_readdata;    // JTAG:av_readdata -> mm_interconnect_0:JTAG_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_avalon_jtag_slave_waitrequest; // JTAG:av_waitrequest -> mm_interconnect_0:JTAG_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_avalon_jtag_slave_address;     // mm_interconnect_0:JTAG_avalon_jtag_slave_address -> JTAG:av_address
	wire         mm_interconnect_0_jtag_avalon_jtag_slave_read;        // mm_interconnect_0:JTAG_avalon_jtag_slave_read -> JTAG:av_read_n
	wire         mm_interconnect_0_jtag_avalon_jtag_slave_write;       // mm_interconnect_0:JTAG_avalon_jtag_slave_write -> JTAG:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_avalon_jtag_slave_writedata;   // mm_interconnect_0:JTAG_avalon_jtag_slave_writedata -> JTAG:av_writedata
	wire  [31:0] mm_interconnect_0_cpu_debug_mem_slave_readdata;       // CPU:debug_mem_slave_readdata -> mm_interconnect_0:CPU_debug_mem_slave_readdata
	wire         mm_interconnect_0_cpu_debug_mem_slave_waitrequest;    // CPU:debug_mem_slave_waitrequest -> mm_interconnect_0:CPU_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_cpu_debug_mem_slave_debugaccess;    // mm_interconnect_0:CPU_debug_mem_slave_debugaccess -> CPU:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_cpu_debug_mem_slave_address;        // mm_interconnect_0:CPU_debug_mem_slave_address -> CPU:debug_mem_slave_address
	wire         mm_interconnect_0_cpu_debug_mem_slave_read;           // mm_interconnect_0:CPU_debug_mem_slave_read -> CPU:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_cpu_debug_mem_slave_byteenable;     // mm_interconnect_0:CPU_debug_mem_slave_byteenable -> CPU:debug_mem_slave_byteenable
	wire         mm_interconnect_0_cpu_debug_mem_slave_write;          // mm_interconnect_0:CPU_debug_mem_slave_write -> CPU:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_cpu_debug_mem_slave_writedata;      // mm_interconnect_0:CPU_debug_mem_slave_writedata -> CPU:debug_mem_slave_writedata
	wire         mm_interconnect_0_ram_s1_chipselect;                  // mm_interconnect_0:RAM_s1_chipselect -> RAM:chipselect
	wire  [31:0] mm_interconnect_0_ram_s1_readdata;                    // RAM:readdata -> mm_interconnect_0:RAM_s1_readdata
	wire  [11:0] mm_interconnect_0_ram_s1_address;                     // mm_interconnect_0:RAM_s1_address -> RAM:address
	wire   [3:0] mm_interconnect_0_ram_s1_byteenable;                  // mm_interconnect_0:RAM_s1_byteenable -> RAM:byteenable
	wire         mm_interconnect_0_ram_s1_write;                       // mm_interconnect_0:RAM_s1_write -> RAM:write
	wire  [31:0] mm_interconnect_0_ram_s1_writedata;                   // mm_interconnect_0:RAM_s1_writedata -> RAM:writedata
	wire         mm_interconnect_0_ram_s1_clken;                       // mm_interconnect_0:RAM_s1_clken -> RAM:clken
	wire         mm_interconnect_0_seg_1_s1_chipselect;                // mm_interconnect_0:SEG_1_s1_chipselect -> SEG_1:chipselect
	wire  [31:0] mm_interconnect_0_seg_1_s1_readdata;                  // SEG_1:readdata -> mm_interconnect_0:SEG_1_s1_readdata
	wire   [1:0] mm_interconnect_0_seg_1_s1_address;                   // mm_interconnect_0:SEG_1_s1_address -> SEG_1:address
	wire         mm_interconnect_0_seg_1_s1_write;                     // mm_interconnect_0:SEG_1_s1_write -> SEG_1:write_n
	wire  [31:0] mm_interconnect_0_seg_1_s1_writedata;                 // mm_interconnect_0:SEG_1_s1_writedata -> SEG_1:writedata
	wire         mm_interconnect_0_timer_s1_chipselect;                // mm_interconnect_0:Timer_s1_chipselect -> Timer:chipselect
	wire  [15:0] mm_interconnect_0_timer_s1_readdata;                  // Timer:readdata -> mm_interconnect_0:Timer_s1_readdata
	wire   [2:0] mm_interconnect_0_timer_s1_address;                   // mm_interconnect_0:Timer_s1_address -> Timer:address
	wire         mm_interconnect_0_timer_s1_write;                     // mm_interconnect_0:Timer_s1_write -> Timer:write_n
	wire  [15:0] mm_interconnect_0_timer_s1_writedata;                 // mm_interconnect_0:Timer_s1_writedata -> Timer:writedata
	wire         mm_interconnect_0_seg_2_s1_chipselect;                // mm_interconnect_0:SEG_2_s1_chipselect -> SEG_2:chipselect
	wire  [31:0] mm_interconnect_0_seg_2_s1_readdata;                  // SEG_2:readdata -> mm_interconnect_0:SEG_2_s1_readdata
	wire   [1:0] mm_interconnect_0_seg_2_s1_address;                   // mm_interconnect_0:SEG_2_s1_address -> SEG_2:address
	wire         mm_interconnect_0_seg_2_s1_write;                     // mm_interconnect_0:SEG_2_s1_write -> SEG_2:write_n
	wire  [31:0] mm_interconnect_0_seg_2_s1_writedata;                 // mm_interconnect_0:SEG_2_s1_writedata -> SEG_2:writedata
	wire         mm_interconnect_0_seg_3_s1_chipselect;                // mm_interconnect_0:SEG_3_s1_chipselect -> SEG_3:chipselect
	wire  [31:0] mm_interconnect_0_seg_3_s1_readdata;                  // SEG_3:readdata -> mm_interconnect_0:SEG_3_s1_readdata
	wire   [1:0] mm_interconnect_0_seg_3_s1_address;                   // mm_interconnect_0:SEG_3_s1_address -> SEG_3:address
	wire         mm_interconnect_0_seg_3_s1_write;                     // mm_interconnect_0:SEG_3_s1_write -> SEG_3:write_n
	wire  [31:0] mm_interconnect_0_seg_3_s1_writedata;                 // mm_interconnect_0:SEG_3_s1_writedata -> SEG_3:writedata
	wire         mm_interconnect_0_seg_4_s1_chipselect;                // mm_interconnect_0:SEG_4_s1_chipselect -> SEG_4:chipselect
	wire  [31:0] mm_interconnect_0_seg_4_s1_readdata;                  // SEG_4:readdata -> mm_interconnect_0:SEG_4_s1_readdata
	wire   [1:0] mm_interconnect_0_seg_4_s1_address;                   // mm_interconnect_0:SEG_4_s1_address -> SEG_4:address
	wire         mm_interconnect_0_seg_4_s1_write;                     // mm_interconnect_0:SEG_4_s1_write -> SEG_4:write_n
	wire  [31:0] mm_interconnect_0_seg_4_s1_writedata;                 // mm_interconnect_0:SEG_4_s1_writedata -> SEG_4:writedata
	wire         mm_interconnect_0_seg_5_s1_chipselect;                // mm_interconnect_0:SEG_5_s1_chipselect -> SEG_5:chipselect
	wire  [31:0] mm_interconnect_0_seg_5_s1_readdata;                  // SEG_5:readdata -> mm_interconnect_0:SEG_5_s1_readdata
	wire   [1:0] mm_interconnect_0_seg_5_s1_address;                   // mm_interconnect_0:SEG_5_s1_address -> SEG_5:address
	wire         mm_interconnect_0_seg_5_s1_write;                     // mm_interconnect_0:SEG_5_s1_write -> SEG_5:write_n
	wire  [31:0] mm_interconnect_0_seg_5_s1_writedata;                 // mm_interconnect_0:SEG_5_s1_writedata -> SEG_5:writedata
	wire         mm_interconnect_0_seg_6_s1_chipselect;                // mm_interconnect_0:SEG_6_s1_chipselect -> SEG_6:chipselect
	wire  [31:0] mm_interconnect_0_seg_6_s1_readdata;                  // SEG_6:readdata -> mm_interconnect_0:SEG_6_s1_readdata
	wire   [1:0] mm_interconnect_0_seg_6_s1_address;                   // mm_interconnect_0:SEG_6_s1_address -> SEG_6:address
	wire         mm_interconnect_0_seg_6_s1_write;                     // mm_interconnect_0:SEG_6_s1_write -> SEG_6:write_n
	wire  [31:0] mm_interconnect_0_seg_6_s1_writedata;                 // mm_interconnect_0:SEG_6_s1_writedata -> SEG_6:writedata
	wire         mm_interconnect_0_leds_s1_chipselect;                 // mm_interconnect_0:LEDS_s1_chipselect -> LEDS:chipselect
	wire  [31:0] mm_interconnect_0_leds_s1_readdata;                   // LEDS:readdata -> mm_interconnect_0:LEDS_s1_readdata
	wire   [1:0] mm_interconnect_0_leds_s1_address;                    // mm_interconnect_0:LEDS_s1_address -> LEDS:address
	wire         mm_interconnect_0_leds_s1_write;                      // mm_interconnect_0:LEDS_s1_write -> LEDS:write_n
	wire  [31:0] mm_interconnect_0_leds_s1_writedata;                  // mm_interconnect_0:LEDS_s1_writedata -> LEDS:writedata
	wire         mm_interconnect_0_piorightbutton_s1_chipselect;       // mm_interconnect_0:PioRightButton_s1_chipselect -> PioRightButton:chipselect
	wire  [31:0] mm_interconnect_0_piorightbutton_s1_readdata;         // PioRightButton:readdata -> mm_interconnect_0:PioRightButton_s1_readdata
	wire   [1:0] mm_interconnect_0_piorightbutton_s1_address;          // mm_interconnect_0:PioRightButton_s1_address -> PioRightButton:address
	wire         mm_interconnect_0_piorightbutton_s1_write;            // mm_interconnect_0:PioRightButton_s1_write -> PioRightButton:write_n
	wire  [31:0] mm_interconnect_0_piorightbutton_s1_writedata;        // mm_interconnect_0:PioRightButton_s1_writedata -> PioRightButton:writedata
	wire         mm_interconnect_0_pioupbutton_s1_chipselect;          // mm_interconnect_0:PioUpButton_s1_chipselect -> PioUpButton:chipselect
	wire  [31:0] mm_interconnect_0_pioupbutton_s1_readdata;            // PioUpButton:readdata -> mm_interconnect_0:PioUpButton_s1_readdata
	wire   [1:0] mm_interconnect_0_pioupbutton_s1_address;             // mm_interconnect_0:PioUpButton_s1_address -> PioUpButton:address
	wire         mm_interconnect_0_pioupbutton_s1_write;               // mm_interconnect_0:PioUpButton_s1_write -> PioUpButton:write_n
	wire  [31:0] mm_interconnect_0_pioupbutton_s1_writedata;           // mm_interconnect_0:PioUpButton_s1_writedata -> PioUpButton:writedata
	wire         mm_interconnect_0_piodownbutton_s1_chipselect;        // mm_interconnect_0:PioDownButton_s1_chipselect -> PioDownButton:chipselect
	wire  [31:0] mm_interconnect_0_piodownbutton_s1_readdata;          // PioDownButton:readdata -> mm_interconnect_0:PioDownButton_s1_readdata
	wire   [1:0] mm_interconnect_0_piodownbutton_s1_address;           // mm_interconnect_0:PioDownButton_s1_address -> PioDownButton:address
	wire         mm_interconnect_0_piodownbutton_s1_write;             // mm_interconnect_0:PioDownButton_s1_write -> PioDownButton:write_n
	wire  [31:0] mm_interconnect_0_piodownbutton_s1_writedata;         // mm_interconnect_0:PioDownButton_s1_writedata -> PioDownButton:writedata
	wire         mm_interconnect_0_alarmactiveswitch_s1_chipselect;    // mm_interconnect_0:AlarmActiveSwitch_s1_chipselect -> AlarmActiveSwitch:chipselect
	wire  [31:0] mm_interconnect_0_alarmactiveswitch_s1_readdata;      // AlarmActiveSwitch:readdata -> mm_interconnect_0:AlarmActiveSwitch_s1_readdata
	wire   [1:0] mm_interconnect_0_alarmactiveswitch_s1_address;       // mm_interconnect_0:AlarmActiveSwitch_s1_address -> AlarmActiveSwitch:address
	wire         mm_interconnect_0_alarmactiveswitch_s1_write;         // mm_interconnect_0:AlarmActiveSwitch_s1_write -> AlarmActiveSwitch:write_n
	wire  [31:0] mm_interconnect_0_alarmactiveswitch_s1_writedata;     // mm_interconnect_0:AlarmActiveSwitch_s1_writedata -> AlarmActiveSwitch:writedata
	wire         mm_interconnect_0_timeractiveswitch_s1_chipselect;    // mm_interconnect_0:TimerActiveSwitch_s1_chipselect -> TimerActiveSwitch:chipselect
	wire  [31:0] mm_interconnect_0_timeractiveswitch_s1_readdata;      // TimerActiveSwitch:readdata -> mm_interconnect_0:TimerActiveSwitch_s1_readdata
	wire   [1:0] mm_interconnect_0_timeractiveswitch_s1_address;       // mm_interconnect_0:TimerActiveSwitch_s1_address -> TimerActiveSwitch:address
	wire         mm_interconnect_0_timeractiveswitch_s1_write;         // mm_interconnect_0:TimerActiveSwitch_s1_write -> TimerActiveSwitch:write_n
	wire  [31:0] mm_interconnect_0_timeractiveswitch_s1_writedata;     // mm_interconnect_0:TimerActiveSwitch_s1_writedata -> TimerActiveSwitch:writedata
	wire         mm_interconnect_0_editalarmswitch_s1_chipselect;      // mm_interconnect_0:EditAlarmSwitch_s1_chipselect -> EditAlarmSwitch:chipselect
	wire  [31:0] mm_interconnect_0_editalarmswitch_s1_readdata;        // EditAlarmSwitch:readdata -> mm_interconnect_0:EditAlarmSwitch_s1_readdata
	wire   [1:0] mm_interconnect_0_editalarmswitch_s1_address;         // mm_interconnect_0:EditAlarmSwitch_s1_address -> EditAlarmSwitch:address
	wire         mm_interconnect_0_editalarmswitch_s1_write;           // mm_interconnect_0:EditAlarmSwitch_s1_write -> EditAlarmSwitch:write_n
	wire  [31:0] mm_interconnect_0_editalarmswitch_s1_writedata;       // mm_interconnect_0:EditAlarmSwitch_s1_writedata -> EditAlarmSwitch:writedata
	wire         mm_interconnect_0_pioleftbutton_s1_chipselect;        // mm_interconnect_0:PioLeftButton_s1_chipselect -> PioLeftButton:chipselect
	wire  [31:0] mm_interconnect_0_pioleftbutton_s1_readdata;          // PioLeftButton:readdata -> mm_interconnect_0:PioLeftButton_s1_readdata
	wire   [1:0] mm_interconnect_0_pioleftbutton_s1_address;           // mm_interconnect_0:PioLeftButton_s1_address -> PioLeftButton:address
	wire         mm_interconnect_0_pioleftbutton_s1_write;             // mm_interconnect_0:PioLeftButton_s1_write -> PioLeftButton:write_n
	wire  [31:0] mm_interconnect_0_pioleftbutton_s1_writedata;         // mm_interconnect_0:PioLeftButton_s1_writedata -> PioLeftButton:writedata
	wire         mm_interconnect_0_edittimerswitch_s1_chipselect;      // mm_interconnect_0:EditTimerSwitch_s1_chipselect -> EditTimerSwitch:chipselect
	wire  [31:0] mm_interconnect_0_edittimerswitch_s1_readdata;        // EditTimerSwitch:readdata -> mm_interconnect_0:EditTimerSwitch_s1_readdata
	wire   [1:0] mm_interconnect_0_edittimerswitch_s1_address;         // mm_interconnect_0:EditTimerSwitch_s1_address -> EditTimerSwitch:address
	wire         mm_interconnect_0_edittimerswitch_s1_write;           // mm_interconnect_0:EditTimerSwitch_s1_write -> EditTimerSwitch:write_n
	wire  [31:0] mm_interconnect_0_edittimerswitch_s1_writedata;       // mm_interconnect_0:EditTimerSwitch_s1_writedata -> EditTimerSwitch:writedata
	wire         mm_interconnect_0_edittimeswitch_s1_chipselect;       // mm_interconnect_0:EditTimeSwitch_s1_chipselect -> EditTimeSwitch:chipselect
	wire  [31:0] mm_interconnect_0_edittimeswitch_s1_readdata;         // EditTimeSwitch:readdata -> mm_interconnect_0:EditTimeSwitch_s1_readdata
	wire   [1:0] mm_interconnect_0_edittimeswitch_s1_address;          // mm_interconnect_0:EditTimeSwitch_s1_address -> EditTimeSwitch:address
	wire         mm_interconnect_0_edittimeswitch_s1_write;            // mm_interconnect_0:EditTimeSwitch_s1_write -> EditTimeSwitch:write_n
	wire  [31:0] mm_interconnect_0_edittimeswitch_s1_writedata;        // mm_interconnect_0:EditTimeSwitch_s1_writedata -> EditTimeSwitch:writedata
	wire         mm_interconnect_0_saveswitch_s1_chipselect;           // mm_interconnect_0:SaveSwitch_s1_chipselect -> SaveSwitch:chipselect
	wire  [31:0] mm_interconnect_0_saveswitch_s1_readdata;             // SaveSwitch:readdata -> mm_interconnect_0:SaveSwitch_s1_readdata
	wire   [1:0] mm_interconnect_0_saveswitch_s1_address;              // mm_interconnect_0:SaveSwitch_s1_address -> SaveSwitch:address
	wire         mm_interconnect_0_saveswitch_s1_write;                // mm_interconnect_0:SaveSwitch_s1_write -> SaveSwitch:write_n
	wire  [31:0] mm_interconnect_0_saveswitch_s1_writedata;            // mm_interconnect_0:SaveSwitch_s1_writedata -> SaveSwitch:writedata
	wire         mm_interconnect_0_uart_s1_chipselect;                 // mm_interconnect_0:UART_s1_chipselect -> UART:chipselect
	wire  [15:0] mm_interconnect_0_uart_s1_readdata;                   // UART:readdata -> mm_interconnect_0:UART_s1_readdata
	wire   [2:0] mm_interconnect_0_uart_s1_address;                    // mm_interconnect_0:UART_s1_address -> UART:address
	wire         mm_interconnect_0_uart_s1_read;                       // mm_interconnect_0:UART_s1_read -> UART:read_n
	wire         mm_interconnect_0_uart_s1_begintransfer;              // mm_interconnect_0:UART_s1_begintransfer -> UART:begintransfer
	wire         mm_interconnect_0_uart_s1_write;                      // mm_interconnect_0:UART_s1_write -> UART:write_n
	wire  [15:0] mm_interconnect_0_uart_s1_writedata;                  // mm_interconnect_0:UART_s1_writedata -> UART:writedata
	wire         irq_mapper_receiver0_irq;                             // JTAG:av_irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                             // Timer:irq -> irq_mapper:receiver1_irq
	wire         irq_mapper_receiver2_irq;                             // PioRightButton:irq -> irq_mapper:receiver2_irq
	wire         irq_mapper_receiver3_irq;                             // PioUpButton:irq -> irq_mapper:receiver3_irq
	wire         irq_mapper_receiver4_irq;                             // PioDownButton:irq -> irq_mapper:receiver4_irq
	wire         irq_mapper_receiver5_irq;                             // AlarmActiveSwitch:irq -> irq_mapper:receiver5_irq
	wire         irq_mapper_receiver6_irq;                             // TimerActiveSwitch:irq -> irq_mapper:receiver6_irq
	wire         irq_mapper_receiver7_irq;                             // EditAlarmSwitch:irq -> irq_mapper:receiver7_irq
	wire         irq_mapper_receiver8_irq;                             // PioLeftButton:irq -> irq_mapper:receiver8_irq
	wire         irq_mapper_receiver9_irq;                             // EditTimerSwitch:irq -> irq_mapper:receiver9_irq
	wire         irq_mapper_receiver10_irq;                            // EditTimeSwitch:irq -> irq_mapper:receiver10_irq
	wire         irq_mapper_receiver11_irq;                            // SaveSwitch:irq -> irq_mapper:receiver11_irq
	wire         irq_mapper_receiver12_irq;                            // UART:irq -> irq_mapper:receiver12_irq
	wire  [31:0] cpu_irq_irq;                                          // irq_mapper:sender_irq -> CPU:irq
	wire         rst_controller_reset_out_reset;                       // rst_controller:reset_out -> [AlarmActiveSwitch:reset_n, CPU:reset_n, EditAlarmSwitch:reset_n, EditTimeSwitch:reset_n, EditTimerSwitch:reset_n, JTAG:rst_n, LEDS:reset_n, PioDownButton:reset_n, PioLeftButton:reset_n, PioRightButton:reset_n, PioUpButton:reset_n, RAM:reset, SEG_1:reset_n, SEG_2:reset_n, SEG_3:reset_n, SEG_4:reset_n, SEG_5:reset_n, SEG_6:reset_n, SaveSwitch:reset_n, Timer:reset_n, TimerActiveSwitch:reset_n, UART:reset_n, irq_mapper:reset, mm_interconnect_0:CPU_reset_reset_bridge_in_reset_reset, rst_translator:in_reset]
	wire         rst_controller_reset_out_reset_req;                   // rst_controller:reset_req -> [CPU:reset_req, RAM:reset_req, rst_translator:reset_req_in]

	ProjectFile_AlarmActiveSwitch alarmactiveswitch (
		.clk        (clk_clk),                                           //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                   //               reset.reset_n
		.address    (mm_interconnect_0_alarmactiveswitch_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_alarmactiveswitch_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_alarmactiveswitch_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_alarmactiveswitch_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_alarmactiveswitch_s1_readdata),   //                    .readdata
		.in_port    (alarm_active_switch_export),                        // external_connection.export
		.irq        (irq_mapper_receiver5_irq)                           //                 irq.irq
	);

	ProjectFile_CPU cpu (
		.clk                                 (clk_clk),                                           //                       clk.clk
		.reset_n                             (~rst_controller_reset_out_reset),                   //                     reset.reset_n
		.reset_req                           (rst_controller_reset_out_reset_req),                //                          .reset_req
		.d_address                           (cpu_data_master_address),                           //               data_master.address
		.d_byteenable                        (cpu_data_master_byteenable),                        //                          .byteenable
		.d_read                              (cpu_data_master_read),                              //                          .read
		.d_readdata                          (cpu_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (cpu_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (cpu_data_master_write),                             //                          .write
		.d_writedata                         (cpu_data_master_writedata),                         //                          .writedata
		.debug_mem_slave_debugaccess_to_roms (cpu_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (cpu_instruction_master_address),                    //        instruction_master.address
		.i_read                              (cpu_instruction_master_read),                       //                          .read
		.i_readdata                          (cpu_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (cpu_instruction_master_waitrequest),                //                          .waitrequest
		.irq                                 (cpu_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (),                                                  //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_cpu_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_cpu_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_cpu_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_cpu_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_cpu_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_cpu_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_cpu_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_cpu_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                   // custom_instruction_master.readra
	);

	ProjectFile_AlarmActiveSwitch editalarmswitch (
		.clk        (clk_clk),                                         //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                 //               reset.reset_n
		.address    (mm_interconnect_0_editalarmswitch_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_editalarmswitch_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_editalarmswitch_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_editalarmswitch_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_editalarmswitch_s1_readdata),   //                    .readdata
		.in_port    (edit_alarm_switch_export),                        // external_connection.export
		.irq        (irq_mapper_receiver7_irq)                         //                 irq.irq
	);

	ProjectFile_AlarmActiveSwitch edittimeswitch (
		.clk        (clk_clk),                                        //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                //               reset.reset_n
		.address    (mm_interconnect_0_edittimeswitch_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_edittimeswitch_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_edittimeswitch_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_edittimeswitch_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_edittimeswitch_s1_readdata),   //                    .readdata
		.in_port    (edit_time_switch_export),                        // external_connection.export
		.irq        (irq_mapper_receiver10_irq)                       //                 irq.irq
	);

	ProjectFile_AlarmActiveSwitch edittimerswitch (
		.clk        (clk_clk),                                         //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                 //               reset.reset_n
		.address    (mm_interconnect_0_edittimerswitch_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_edittimerswitch_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_edittimerswitch_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_edittimerswitch_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_edittimerswitch_s1_readdata),   //                    .readdata
		.in_port    (edit_timer_switch_export),                        // external_connection.export
		.irq        (irq_mapper_receiver9_irq)                         //                 irq.irq
	);

	ProjectFile_JTAG jtag (
		.clk            (clk_clk),                                              //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                      //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                              //               irq.irq
	);

	ProjectFile_LEDS leds (
		.clk        (clk_clk),                              //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_leds_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_leds_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_leds_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_leds_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_leds_s1_readdata),   //                    .readdata
		.out_port   (leds_export)                           // external_connection.export
	);

	ProjectFile_AlarmActiveSwitch piodownbutton (
		.clk        (clk_clk),                                       //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),               //               reset.reset_n
		.address    (mm_interconnect_0_piodownbutton_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_piodownbutton_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_piodownbutton_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_piodownbutton_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_piodownbutton_s1_readdata),   //                    .readdata
		.in_port    (down_button_export),                            // external_connection.export
		.irq        (irq_mapper_receiver4_irq)                       //                 irq.irq
	);

	ProjectFile_AlarmActiveSwitch pioleftbutton (
		.clk        (clk_clk),                                       //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),               //               reset.reset_n
		.address    (mm_interconnect_0_pioleftbutton_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_pioleftbutton_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_pioleftbutton_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_pioleftbutton_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_pioleftbutton_s1_readdata),   //                    .readdata
		.in_port    (left_button_export),                            // external_connection.export
		.irq        (irq_mapper_receiver8_irq)                       //                 irq.irq
	);

	ProjectFile_AlarmActiveSwitch piorightbutton (
		.clk        (clk_clk),                                        //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                //               reset.reset_n
		.address    (mm_interconnect_0_piorightbutton_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_piorightbutton_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_piorightbutton_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_piorightbutton_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_piorightbutton_s1_readdata),   //                    .readdata
		.in_port    (right_button_export),                            // external_connection.export
		.irq        (irq_mapper_receiver2_irq)                        //                 irq.irq
	);

	ProjectFile_AlarmActiveSwitch pioupbutton (
		.clk        (clk_clk),                                     //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),             //               reset.reset_n
		.address    (mm_interconnect_0_pioupbutton_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_pioupbutton_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_pioupbutton_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_pioupbutton_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_pioupbutton_s1_readdata),   //                    .readdata
		.in_port    (up_button_export),                            // external_connection.export
		.irq        (irq_mapper_receiver3_irq)                     //                 irq.irq
	);

	ProjectFile_RAM ram (
		.clk        (clk_clk),                             //   clk1.clk
		.address    (mm_interconnect_0_ram_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_ram_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_ram_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_ram_s1_write),      //       .write
		.readdata   (mm_interconnect_0_ram_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_ram_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_ram_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),      // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req),  //       .reset_req
		.freeze     (1'b0)                                 // (terminated)
	);

	ProjectFile_SEG_1 seg_1 (
		.clk        (clk_clk),                               //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),       //               reset.reset_n
		.address    (mm_interconnect_0_seg_1_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_seg_1_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_seg_1_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_seg_1_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_seg_1_s1_readdata),   //                    .readdata
		.out_port   (segment1_export)                        // external_connection.export
	);

	ProjectFile_SEG_1 seg_2 (
		.clk        (clk_clk),                               //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),       //               reset.reset_n
		.address    (mm_interconnect_0_seg_2_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_seg_2_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_seg_2_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_seg_2_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_seg_2_s1_readdata),   //                    .readdata
		.out_port   (segment2_export)                        // external_connection.export
	);

	ProjectFile_SEG_1 seg_3 (
		.clk        (clk_clk),                               //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),       //               reset.reset_n
		.address    (mm_interconnect_0_seg_3_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_seg_3_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_seg_3_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_seg_3_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_seg_3_s1_readdata),   //                    .readdata
		.out_port   (segment3_export)                        // external_connection.export
	);

	ProjectFile_SEG_1 seg_4 (
		.clk        (clk_clk),                               //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),       //               reset.reset_n
		.address    (mm_interconnect_0_seg_4_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_seg_4_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_seg_4_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_seg_4_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_seg_4_s1_readdata),   //                    .readdata
		.out_port   (segment4_export)                        // external_connection.export
	);

	ProjectFile_SEG_1 seg_5 (
		.clk        (clk_clk),                               //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),       //               reset.reset_n
		.address    (mm_interconnect_0_seg_5_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_seg_5_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_seg_5_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_seg_5_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_seg_5_s1_readdata),   //                    .readdata
		.out_port   (segment5_export)                        // external_connection.export
	);

	ProjectFile_SEG_1 seg_6 (
		.clk        (clk_clk),                               //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),       //               reset.reset_n
		.address    (mm_interconnect_0_seg_6_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_seg_6_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_seg_6_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_seg_6_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_seg_6_s1_readdata),   //                    .readdata
		.out_port   (segment6_export)                        // external_connection.export
	);

	ProjectFile_AlarmActiveSwitch saveswitch (
		.clk        (clk_clk),                                    //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),            //               reset.reset_n
		.address    (mm_interconnect_0_saveswitch_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_saveswitch_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_saveswitch_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_saveswitch_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_saveswitch_s1_readdata),   //                    .readdata
		.in_port    (save_switch_export),                         // external_connection.export
		.irq        (irq_mapper_receiver11_irq)                   //                 irq.irq
	);

	ProjectFile_Timer timer (
		.clk        (clk_clk),                               //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),       // reset.reset_n
		.address    (mm_interconnect_0_timer_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timer_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timer_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timer_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timer_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver1_irq)               //   irq.irq
	);

	ProjectFile_AlarmActiveSwitch timeractiveswitch (
		.clk        (clk_clk),                                           //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                   //               reset.reset_n
		.address    (mm_interconnect_0_timeractiveswitch_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_timeractiveswitch_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_timeractiveswitch_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_timeractiveswitch_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_timeractiveswitch_s1_readdata),   //                    .readdata
		.in_port    (timer_active_switch_export),                        // external_connection.export
		.irq        (irq_mapper_receiver6_irq)                           //                 irq.irq
	);

	ProjectFile_UART uart (
		.clk           (clk_clk),                                 //                 clk.clk
		.reset_n       (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address       (mm_interconnect_0_uart_s1_address),       //                  s1.address
		.begintransfer (mm_interconnect_0_uart_s1_begintransfer), //                    .begintransfer
		.chipselect    (mm_interconnect_0_uart_s1_chipselect),    //                    .chipselect
		.read_n        (~mm_interconnect_0_uart_s1_read),         //                    .read_n
		.write_n       (~mm_interconnect_0_uart_s1_write),        //                    .write_n
		.writedata     (mm_interconnect_0_uart_s1_writedata),     //                    .writedata
		.readdata      (mm_interconnect_0_uart_s1_readdata),      //                    .readdata
		.rxd           (uart_rxd),                                // external_connection.export
		.txd           (uart_txd),                                //                    .export
		.irq           (irq_mapper_receiver12_irq)                //                 irq.irq
	);

	ProjectFile_mm_interconnect_0 mm_interconnect_0 (
		.CLK_clk_clk                           (clk_clk),                                              //                         CLK_clk.clk
		.CPU_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                       // CPU_reset_reset_bridge_in_reset.reset
		.CPU_data_master_address               (cpu_data_master_address),                              //                 CPU_data_master.address
		.CPU_data_master_waitrequest           (cpu_data_master_waitrequest),                          //                                .waitrequest
		.CPU_data_master_byteenable            (cpu_data_master_byteenable),                           //                                .byteenable
		.CPU_data_master_read                  (cpu_data_master_read),                                 //                                .read
		.CPU_data_master_readdata              (cpu_data_master_readdata),                             //                                .readdata
		.CPU_data_master_write                 (cpu_data_master_write),                                //                                .write
		.CPU_data_master_writedata             (cpu_data_master_writedata),                            //                                .writedata
		.CPU_data_master_debugaccess           (cpu_data_master_debugaccess),                          //                                .debugaccess
		.CPU_instruction_master_address        (cpu_instruction_master_address),                       //          CPU_instruction_master.address
		.CPU_instruction_master_waitrequest    (cpu_instruction_master_waitrequest),                   //                                .waitrequest
		.CPU_instruction_master_read           (cpu_instruction_master_read),                          //                                .read
		.CPU_instruction_master_readdata       (cpu_instruction_master_readdata),                      //                                .readdata
		.AlarmActiveSwitch_s1_address          (mm_interconnect_0_alarmactiveswitch_s1_address),       //            AlarmActiveSwitch_s1.address
		.AlarmActiveSwitch_s1_write            (mm_interconnect_0_alarmactiveswitch_s1_write),         //                                .write
		.AlarmActiveSwitch_s1_readdata         (mm_interconnect_0_alarmactiveswitch_s1_readdata),      //                                .readdata
		.AlarmActiveSwitch_s1_writedata        (mm_interconnect_0_alarmactiveswitch_s1_writedata),     //                                .writedata
		.AlarmActiveSwitch_s1_chipselect       (mm_interconnect_0_alarmactiveswitch_s1_chipselect),    //                                .chipselect
		.CPU_debug_mem_slave_address           (mm_interconnect_0_cpu_debug_mem_slave_address),        //             CPU_debug_mem_slave.address
		.CPU_debug_mem_slave_write             (mm_interconnect_0_cpu_debug_mem_slave_write),          //                                .write
		.CPU_debug_mem_slave_read              (mm_interconnect_0_cpu_debug_mem_slave_read),           //                                .read
		.CPU_debug_mem_slave_readdata          (mm_interconnect_0_cpu_debug_mem_slave_readdata),       //                                .readdata
		.CPU_debug_mem_slave_writedata         (mm_interconnect_0_cpu_debug_mem_slave_writedata),      //                                .writedata
		.CPU_debug_mem_slave_byteenable        (mm_interconnect_0_cpu_debug_mem_slave_byteenable),     //                                .byteenable
		.CPU_debug_mem_slave_waitrequest       (mm_interconnect_0_cpu_debug_mem_slave_waitrequest),    //                                .waitrequest
		.CPU_debug_mem_slave_debugaccess       (mm_interconnect_0_cpu_debug_mem_slave_debugaccess),    //                                .debugaccess
		.EditAlarmSwitch_s1_address            (mm_interconnect_0_editalarmswitch_s1_address),         //              EditAlarmSwitch_s1.address
		.EditAlarmSwitch_s1_write              (mm_interconnect_0_editalarmswitch_s1_write),           //                                .write
		.EditAlarmSwitch_s1_readdata           (mm_interconnect_0_editalarmswitch_s1_readdata),        //                                .readdata
		.EditAlarmSwitch_s1_writedata          (mm_interconnect_0_editalarmswitch_s1_writedata),       //                                .writedata
		.EditAlarmSwitch_s1_chipselect         (mm_interconnect_0_editalarmswitch_s1_chipselect),      //                                .chipselect
		.EditTimerSwitch_s1_address            (mm_interconnect_0_edittimerswitch_s1_address),         //              EditTimerSwitch_s1.address
		.EditTimerSwitch_s1_write              (mm_interconnect_0_edittimerswitch_s1_write),           //                                .write
		.EditTimerSwitch_s1_readdata           (mm_interconnect_0_edittimerswitch_s1_readdata),        //                                .readdata
		.EditTimerSwitch_s1_writedata          (mm_interconnect_0_edittimerswitch_s1_writedata),       //                                .writedata
		.EditTimerSwitch_s1_chipselect         (mm_interconnect_0_edittimerswitch_s1_chipselect),      //                                .chipselect
		.EditTimeSwitch_s1_address             (mm_interconnect_0_edittimeswitch_s1_address),          //               EditTimeSwitch_s1.address
		.EditTimeSwitch_s1_write               (mm_interconnect_0_edittimeswitch_s1_write),            //                                .write
		.EditTimeSwitch_s1_readdata            (mm_interconnect_0_edittimeswitch_s1_readdata),         //                                .readdata
		.EditTimeSwitch_s1_writedata           (mm_interconnect_0_edittimeswitch_s1_writedata),        //                                .writedata
		.EditTimeSwitch_s1_chipselect          (mm_interconnect_0_edittimeswitch_s1_chipselect),       //                                .chipselect
		.JTAG_avalon_jtag_slave_address        (mm_interconnect_0_jtag_avalon_jtag_slave_address),     //          JTAG_avalon_jtag_slave.address
		.JTAG_avalon_jtag_slave_write          (mm_interconnect_0_jtag_avalon_jtag_slave_write),       //                                .write
		.JTAG_avalon_jtag_slave_read           (mm_interconnect_0_jtag_avalon_jtag_slave_read),        //                                .read
		.JTAG_avalon_jtag_slave_readdata       (mm_interconnect_0_jtag_avalon_jtag_slave_readdata),    //                                .readdata
		.JTAG_avalon_jtag_slave_writedata      (mm_interconnect_0_jtag_avalon_jtag_slave_writedata),   //                                .writedata
		.JTAG_avalon_jtag_slave_waitrequest    (mm_interconnect_0_jtag_avalon_jtag_slave_waitrequest), //                                .waitrequest
		.JTAG_avalon_jtag_slave_chipselect     (mm_interconnect_0_jtag_avalon_jtag_slave_chipselect),  //                                .chipselect
		.LEDS_s1_address                       (mm_interconnect_0_leds_s1_address),                    //                         LEDS_s1.address
		.LEDS_s1_write                         (mm_interconnect_0_leds_s1_write),                      //                                .write
		.LEDS_s1_readdata                      (mm_interconnect_0_leds_s1_readdata),                   //                                .readdata
		.LEDS_s1_writedata                     (mm_interconnect_0_leds_s1_writedata),                  //                                .writedata
		.LEDS_s1_chipselect                    (mm_interconnect_0_leds_s1_chipselect),                 //                                .chipselect
		.PioDownButton_s1_address              (mm_interconnect_0_piodownbutton_s1_address),           //                PioDownButton_s1.address
		.PioDownButton_s1_write                (mm_interconnect_0_piodownbutton_s1_write),             //                                .write
		.PioDownButton_s1_readdata             (mm_interconnect_0_piodownbutton_s1_readdata),          //                                .readdata
		.PioDownButton_s1_writedata            (mm_interconnect_0_piodownbutton_s1_writedata),         //                                .writedata
		.PioDownButton_s1_chipselect           (mm_interconnect_0_piodownbutton_s1_chipselect),        //                                .chipselect
		.PioLeftButton_s1_address              (mm_interconnect_0_pioleftbutton_s1_address),           //                PioLeftButton_s1.address
		.PioLeftButton_s1_write                (mm_interconnect_0_pioleftbutton_s1_write),             //                                .write
		.PioLeftButton_s1_readdata             (mm_interconnect_0_pioleftbutton_s1_readdata),          //                                .readdata
		.PioLeftButton_s1_writedata            (mm_interconnect_0_pioleftbutton_s1_writedata),         //                                .writedata
		.PioLeftButton_s1_chipselect           (mm_interconnect_0_pioleftbutton_s1_chipselect),        //                                .chipselect
		.PioRightButton_s1_address             (mm_interconnect_0_piorightbutton_s1_address),          //               PioRightButton_s1.address
		.PioRightButton_s1_write               (mm_interconnect_0_piorightbutton_s1_write),            //                                .write
		.PioRightButton_s1_readdata            (mm_interconnect_0_piorightbutton_s1_readdata),         //                                .readdata
		.PioRightButton_s1_writedata           (mm_interconnect_0_piorightbutton_s1_writedata),        //                                .writedata
		.PioRightButton_s1_chipselect          (mm_interconnect_0_piorightbutton_s1_chipselect),       //                                .chipselect
		.PioUpButton_s1_address                (mm_interconnect_0_pioupbutton_s1_address),             //                  PioUpButton_s1.address
		.PioUpButton_s1_write                  (mm_interconnect_0_pioupbutton_s1_write),               //                                .write
		.PioUpButton_s1_readdata               (mm_interconnect_0_pioupbutton_s1_readdata),            //                                .readdata
		.PioUpButton_s1_writedata              (mm_interconnect_0_pioupbutton_s1_writedata),           //                                .writedata
		.PioUpButton_s1_chipselect             (mm_interconnect_0_pioupbutton_s1_chipselect),          //                                .chipselect
		.RAM_s1_address                        (mm_interconnect_0_ram_s1_address),                     //                          RAM_s1.address
		.RAM_s1_write                          (mm_interconnect_0_ram_s1_write),                       //                                .write
		.RAM_s1_readdata                       (mm_interconnect_0_ram_s1_readdata),                    //                                .readdata
		.RAM_s1_writedata                      (mm_interconnect_0_ram_s1_writedata),                   //                                .writedata
		.RAM_s1_byteenable                     (mm_interconnect_0_ram_s1_byteenable),                  //                                .byteenable
		.RAM_s1_chipselect                     (mm_interconnect_0_ram_s1_chipselect),                  //                                .chipselect
		.RAM_s1_clken                          (mm_interconnect_0_ram_s1_clken),                       //                                .clken
		.SaveSwitch_s1_address                 (mm_interconnect_0_saveswitch_s1_address),              //                   SaveSwitch_s1.address
		.SaveSwitch_s1_write                   (mm_interconnect_0_saveswitch_s1_write),                //                                .write
		.SaveSwitch_s1_readdata                (mm_interconnect_0_saveswitch_s1_readdata),             //                                .readdata
		.SaveSwitch_s1_writedata               (mm_interconnect_0_saveswitch_s1_writedata),            //                                .writedata
		.SaveSwitch_s1_chipselect              (mm_interconnect_0_saveswitch_s1_chipselect),           //                                .chipselect
		.SEG_1_s1_address                      (mm_interconnect_0_seg_1_s1_address),                   //                        SEG_1_s1.address
		.SEG_1_s1_write                        (mm_interconnect_0_seg_1_s1_write),                     //                                .write
		.SEG_1_s1_readdata                     (mm_interconnect_0_seg_1_s1_readdata),                  //                                .readdata
		.SEG_1_s1_writedata                    (mm_interconnect_0_seg_1_s1_writedata),                 //                                .writedata
		.SEG_1_s1_chipselect                   (mm_interconnect_0_seg_1_s1_chipselect),                //                                .chipselect
		.SEG_2_s1_address                      (mm_interconnect_0_seg_2_s1_address),                   //                        SEG_2_s1.address
		.SEG_2_s1_write                        (mm_interconnect_0_seg_2_s1_write),                     //                                .write
		.SEG_2_s1_readdata                     (mm_interconnect_0_seg_2_s1_readdata),                  //                                .readdata
		.SEG_2_s1_writedata                    (mm_interconnect_0_seg_2_s1_writedata),                 //                                .writedata
		.SEG_2_s1_chipselect                   (mm_interconnect_0_seg_2_s1_chipselect),                //                                .chipselect
		.SEG_3_s1_address                      (mm_interconnect_0_seg_3_s1_address),                   //                        SEG_3_s1.address
		.SEG_3_s1_write                        (mm_interconnect_0_seg_3_s1_write),                     //                                .write
		.SEG_3_s1_readdata                     (mm_interconnect_0_seg_3_s1_readdata),                  //                                .readdata
		.SEG_3_s1_writedata                    (mm_interconnect_0_seg_3_s1_writedata),                 //                                .writedata
		.SEG_3_s1_chipselect                   (mm_interconnect_0_seg_3_s1_chipselect),                //                                .chipselect
		.SEG_4_s1_address                      (mm_interconnect_0_seg_4_s1_address),                   //                        SEG_4_s1.address
		.SEG_4_s1_write                        (mm_interconnect_0_seg_4_s1_write),                     //                                .write
		.SEG_4_s1_readdata                     (mm_interconnect_0_seg_4_s1_readdata),                  //                                .readdata
		.SEG_4_s1_writedata                    (mm_interconnect_0_seg_4_s1_writedata),                 //                                .writedata
		.SEG_4_s1_chipselect                   (mm_interconnect_0_seg_4_s1_chipselect),                //                                .chipselect
		.SEG_5_s1_address                      (mm_interconnect_0_seg_5_s1_address),                   //                        SEG_5_s1.address
		.SEG_5_s1_write                        (mm_interconnect_0_seg_5_s1_write),                     //                                .write
		.SEG_5_s1_readdata                     (mm_interconnect_0_seg_5_s1_readdata),                  //                                .readdata
		.SEG_5_s1_writedata                    (mm_interconnect_0_seg_5_s1_writedata),                 //                                .writedata
		.SEG_5_s1_chipselect                   (mm_interconnect_0_seg_5_s1_chipselect),                //                                .chipselect
		.SEG_6_s1_address                      (mm_interconnect_0_seg_6_s1_address),                   //                        SEG_6_s1.address
		.SEG_6_s1_write                        (mm_interconnect_0_seg_6_s1_write),                     //                                .write
		.SEG_6_s1_readdata                     (mm_interconnect_0_seg_6_s1_readdata),                  //                                .readdata
		.SEG_6_s1_writedata                    (mm_interconnect_0_seg_6_s1_writedata),                 //                                .writedata
		.SEG_6_s1_chipselect                   (mm_interconnect_0_seg_6_s1_chipselect),                //                                .chipselect
		.Timer_s1_address                      (mm_interconnect_0_timer_s1_address),                   //                        Timer_s1.address
		.Timer_s1_write                        (mm_interconnect_0_timer_s1_write),                     //                                .write
		.Timer_s1_readdata                     (mm_interconnect_0_timer_s1_readdata),                  //                                .readdata
		.Timer_s1_writedata                    (mm_interconnect_0_timer_s1_writedata),                 //                                .writedata
		.Timer_s1_chipselect                   (mm_interconnect_0_timer_s1_chipselect),                //                                .chipselect
		.TimerActiveSwitch_s1_address          (mm_interconnect_0_timeractiveswitch_s1_address),       //            TimerActiveSwitch_s1.address
		.TimerActiveSwitch_s1_write            (mm_interconnect_0_timeractiveswitch_s1_write),         //                                .write
		.TimerActiveSwitch_s1_readdata         (mm_interconnect_0_timeractiveswitch_s1_readdata),      //                                .readdata
		.TimerActiveSwitch_s1_writedata        (mm_interconnect_0_timeractiveswitch_s1_writedata),     //                                .writedata
		.TimerActiveSwitch_s1_chipselect       (mm_interconnect_0_timeractiveswitch_s1_chipselect),    //                                .chipselect
		.UART_s1_address                       (mm_interconnect_0_uart_s1_address),                    //                         UART_s1.address
		.UART_s1_write                         (mm_interconnect_0_uart_s1_write),                      //                                .write
		.UART_s1_read                          (mm_interconnect_0_uart_s1_read),                       //                                .read
		.UART_s1_readdata                      (mm_interconnect_0_uart_s1_readdata),                   //                                .readdata
		.UART_s1_writedata                     (mm_interconnect_0_uart_s1_writedata),                  //                                .writedata
		.UART_s1_begintransfer                 (mm_interconnect_0_uart_s1_begintransfer),              //                                .begintransfer
		.UART_s1_chipselect                    (mm_interconnect_0_uart_s1_chipselect)                  //                                .chipselect
	);

	ProjectFile_irq_mapper irq_mapper (
		.clk            (clk_clk),                        //        clk.clk
		.reset          (rst_controller_reset_out_reset), //  clk_reset.reset
		.receiver0_irq  (irq_mapper_receiver0_irq),       //  receiver0.irq
		.receiver1_irq  (irq_mapper_receiver1_irq),       //  receiver1.irq
		.receiver2_irq  (irq_mapper_receiver2_irq),       //  receiver2.irq
		.receiver3_irq  (irq_mapper_receiver3_irq),       //  receiver3.irq
		.receiver4_irq  (irq_mapper_receiver4_irq),       //  receiver4.irq
		.receiver5_irq  (irq_mapper_receiver5_irq),       //  receiver5.irq
		.receiver6_irq  (irq_mapper_receiver6_irq),       //  receiver6.irq
		.receiver7_irq  (irq_mapper_receiver7_irq),       //  receiver7.irq
		.receiver8_irq  (irq_mapper_receiver8_irq),       //  receiver8.irq
		.receiver9_irq  (irq_mapper_receiver9_irq),       //  receiver9.irq
		.receiver10_irq (irq_mapper_receiver10_irq),      // receiver10.irq
		.receiver11_irq (irq_mapper_receiver11_irq),      // receiver11.irq
		.receiver12_irq (irq_mapper_receiver12_irq),      // receiver12.irq
		.sender_irq     (cpu_irq_irq)                     //     sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
