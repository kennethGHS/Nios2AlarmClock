// ProjectFile_tb.v

// Generated using ACDS version 20.1 720

`timescale 1 ps / 1 ps
module ProjectFile_tb (
	);

	wire        projectfile_inst_clk_bfm_clk_clk;                   // ProjectFile_inst_clk_bfm:clk -> [ProjectFile_inst:clk_clk, ProjectFile_inst_reset_bfm:clk]
	wire  [0:0] projectfile_inst_interrupbutton_bfm_conduit_export; // ProjectFile_inst_interrupbutton_bfm:sig_export -> ProjectFile_inst:interrupbutton_export
	wire  [9:0] projectfile_inst_leds_export;                       // ProjectFile_inst:leds_export -> ProjectFile_inst_leds_bfm:sig_export
	wire  [7:0] projectfile_inst_segment1_export;                   // ProjectFile_inst:segment1_export -> ProjectFile_inst_segment1_bfm:sig_export
	wire  [7:0] projectfile_inst_segment2_export;                   // ProjectFile_inst:segment2_export -> ProjectFile_inst_segment2_bfm:sig_export
	wire  [7:0] projectfile_inst_segment3_export;                   // ProjectFile_inst:segment3_export -> ProjectFile_inst_segment3_bfm:sig_export
	wire  [7:0] projectfile_inst_segment4_export;                   // ProjectFile_inst:segment4_export -> ProjectFile_inst_segment4_bfm:sig_export
	wire  [7:0] projectfile_inst_segment5_export;                   // ProjectFile_inst:segment5_export -> ProjectFile_inst_segment5_bfm:sig_export
	wire  [7:0] projectfile_inst_segment6_export;                   // ProjectFile_inst:segment6_export -> ProjectFile_inst_segment6_bfm:sig_export
	wire        projectfile_inst_uart_txd;                          // ProjectFile_inst:uart_txd -> ProjectFile_inst_uart_bfm:sig_txd
	wire  [0:0] projectfile_inst_uart_bfm_conduit_rxd;              // ProjectFile_inst_uart_bfm:sig_rxd -> ProjectFile_inst:uart_rxd
	wire        projectfile_inst_reset_bfm_reset_reset;             // ProjectFile_inst_reset_bfm:reset -> ProjectFile_inst:reset_reset_n

	ProjectFile projectfile_inst (
		.clk_clk               (projectfile_inst_clk_bfm_clk_clk),                   //            clk.clk
		.interrupbutton_export (projectfile_inst_interrupbutton_bfm_conduit_export), // interrupbutton.export
		.leds_export           (projectfile_inst_leds_export),                       //           leds.export
		.reset_reset_n         (projectfile_inst_reset_bfm_reset_reset),             //          reset.reset_n
		.segment1_export       (projectfile_inst_segment1_export),                   //       segment1.export
		.segment2_export       (projectfile_inst_segment2_export),                   //       segment2.export
		.segment3_export       (projectfile_inst_segment3_export),                   //       segment3.export
		.segment4_export       (projectfile_inst_segment4_export),                   //       segment4.export
		.segment5_export       (projectfile_inst_segment5_export),                   //       segment5.export
		.segment6_export       (projectfile_inst_segment6_export),                   //       segment6.export
		.uart_rxd              (projectfile_inst_uart_bfm_conduit_rxd),              //           uart.rxd
		.uart_txd              (projectfile_inst_uart_txd)                           //               .txd
	);

	altera_avalon_clock_source #(
		.CLOCK_RATE (50000000),
		.CLOCK_UNIT (1)
	) projectfile_inst_clk_bfm (
		.clk (projectfile_inst_clk_bfm_clk_clk)  // clk.clk
	);

	altera_conduit_bfm projectfile_inst_interrupbutton_bfm (
		.sig_export (projectfile_inst_interrupbutton_bfm_conduit_export)  // conduit.export
	);

	altera_conduit_bfm_0002 projectfile_inst_leds_bfm (
		.sig_export (projectfile_inst_leds_export)  // conduit.export
	);

	altera_avalon_reset_source #(
		.ASSERT_HIGH_RESET    (0),
		.INITIAL_RESET_CYCLES (50)
	) projectfile_inst_reset_bfm (
		.reset (projectfile_inst_reset_bfm_reset_reset), // reset.reset_n
		.clk   (projectfile_inst_clk_bfm_clk_clk)        //   clk.clk
	);

	altera_conduit_bfm_0003 projectfile_inst_segment1_bfm (
		.sig_export (projectfile_inst_segment1_export)  // conduit.export
	);

	altera_conduit_bfm_0003 projectfile_inst_segment2_bfm (
		.sig_export (projectfile_inst_segment2_export)  // conduit.export
	);

	altera_conduit_bfm_0003 projectfile_inst_segment3_bfm (
		.sig_export (projectfile_inst_segment3_export)  // conduit.export
	);

	altera_conduit_bfm_0003 projectfile_inst_segment4_bfm (
		.sig_export (projectfile_inst_segment4_export)  // conduit.export
	);

	altera_conduit_bfm_0003 projectfile_inst_segment5_bfm (
		.sig_export (projectfile_inst_segment5_export)  // conduit.export
	);

	altera_conduit_bfm_0003 projectfile_inst_segment6_bfm (
		.sig_export (projectfile_inst_segment6_export)  // conduit.export
	);

	altera_conduit_bfm_0004 projectfile_inst_uart_bfm (
		.sig_rxd (projectfile_inst_uart_bfm_conduit_rxd), // conduit.rxd
		.sig_txd (projectfile_inst_uart_txd)              //        .txd
	);

endmodule
